module top( 
        input   clk,
        input   rstn,
        output  led5,
        output  led6
);
assign led5  =1;
assign led6=0;

endmodule
